//Yarin Digmi 208278655 NIck Garber 322332628
// `timescale  1ns/1ps

module Sum #(
    parameter NOF_BITS = 32
) (
    input wire clk,
    input wire rst_n,
    input wire data_first,
    input wire data_last,
    input wire [NOF_BITS-1:0] data_in,
    output reg [NOF_BITS:0] data_out,
    output reg busy,
    output reg done
);

localparam  READY=0, WORKING=1, FINISH=2;
reg [1:0]state, next_state;
reg [NOF_BITS:0]temp_sum;

always @(*)begin
    data_out={ (NOF_BITS+1){1'b0} };
    done=1'b0;
    busy=1'b0;
    next_state=state;
    case(state)
    READY:begin
        done=1'b0;
        busy=1'b0;
        if(data_first && data_last) next_state=FINISH;
        else if(data_first) next_state=WORKING;
        else next_state=state;
    end
    WORKING:begin
        done=1'b0;
        busy=1'b1;
        if(data_last) next_state=FINISH;
        else next_state=state;
    end
    FINISH:begin
        done=1'b1;
        busy=1'b1;
        next_state=READY;
        data_out= temp_sum;
    end
    endcase
end

always @(posedge clk or negedge rst_n)begin
    if(!rst_n)begin
        state<=READY;
        temp_sum<=0;
    end
    else if(state==READY && data_first)begin
        state<=next_state;
        temp_sum<=data_in;
    end
    else if (state==READY)begin
        state<=next_state;
        temp_sum<=0;
    end
    else begin
        state<=next_state;
        temp_sum<=temp_sum+data_in;
    end
end



endmodule
